a   �	  a   v   F  c  3  @  r  �  �  �  �  �  S  l  x  �  �  �  B	  ^	  j	  �	     v   FileAndType�   F  �{"baseDir":"G:/Game Development/Unity Projects/Core Projects/TirUtilities/Documentation","file":"api/TirUtilities.Vector3Extensions.yml","type":"article","sourceDir":"api/","destinationDir":"api/"}   c  OriginalFileAndType�   3  �{"baseDir":"G:/Game Development/Unity Projects/Core Projects/TirUtilities/Documentation","file":"api/TirUtilities.Vector3Extensions.yml","type":"article","sourceDir":"api/","destinationDir":"api/"}   @  Key2   r  (~/api/TirUtilities.Vector3Extensions.yml   �  LocalPathFromRoot0   �  &api/TirUtilities.Vector3Extensions.yml   �  LinkToFiles	   �     �  
LinkToUids=   S  ,  g  �  �  �    (  ?  p  �  �  �  &  ;   g  1TirUtilities.Vector3Extensions.Invariant(Vector3)3   �  )TirUtilities.Vector3Extensions.Invariant*   �  Global.Vector3(   �  TirUtilities.Vector3Extensions8     .TirUtilities.Vector3Extensions.IsZero(Vector3)   (  TirUtilities   ?  System.Object1   p  'TirUtilities.Vector3Extensions.NotZero*   �  System.Boolean9   �  /TirUtilities.Vector3Extensions.NotZero(Vector3)0   �  &TirUtilities.Vector3Extensions.IsZero*5   &  +TirUtilities.Vector3Extensions.Abs(Vector3)-   S  #TirUtilities.Vector3Extensions.Abs*   l  FileLinkSources   x  {}   �  UidLinkSources   �  {}   �  Uids�  B	  �[{"name":"TirUtilities.Vector3Extensions","file":"api/TirUtilities.Vector3Extensions.yml"},{"name":"TirUtilities.Vector3Extensions.IsZero(Vector3)","file":"api/TirUtilities.Vector3Extensions.yml"},{"name":"TirUtilities.Vector3Extensions.NotZero(Vector3)","file":"api/TirUtilities.Vector3Extensions.yml"},{"name":"TirUtilities.Vector3Extensions.Invariant(Vector3)","file":"api/TirUtilities.Vector3Extensions.yml"},{"name":"TirUtilities.Vector3Extensions.Abs(Vector3)","file":"api/TirUtilities.Vector3Extensions.yml"},{"name":"TirUtilities.Vector3Extensions.IsZero*","file":"api/TirUtilities.Vector3Extensions.yml"},{"name":"TirUtilities.Vector3Extensions.NotZero*","file":"api/TirUtilities.Vector3Extensions.yml"},{"name":"TirUtilities.Vector3Extensions.Invariant*","file":"api/TirUtilities.Vector3Extensions.yml"},{"name":"TirUtilities.Vector3Extensions.Abs*","file":"api/TirUtilities.Vector3Extensions.yml"}]   ^	  ManifestProperties   j	  {}   �	  DocumentType	   �	   �5  s?  {"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.PageViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","items":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"TirUtilities.Vector3Extensions","commentId":"T:TirUtilities.Vector3Extensions","id":"Vector3Extensions","isEii":false,"isExtensionMethod":false,"parent":"TirUtilities","children":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["TirUtilities.Vector3Extensions.Abs(Vector3)","TirUtilities.Vector3Extensions.Invariant(Vector3)","TirUtilities.Vector3Extensions.IsZero(Vector3)","TirUtilities.Vector3Extensions.NotZero(Vector3)"]},"langs":{"$type":"System.String[], mscorlib","$values":["csharp","vb"]},"name":"Vector3Extensions","nameWithType":"Vector3Extensions","fullName":"TirUtilities.Vector3Extensions","type":"Class","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"Vector3Extensions","path":"","startLine":5110,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["cs.temp.dll"]},"namespace":"TirUtilities","summary":"","example":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":[]},"syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public static class Vector3Extensions","content.vb":"Public Module Vector3Extensions"},"inheritance":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["System.Object"]},"modifiers.csharp":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["public","static","class"]},"modifiers.vb":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["Public","Module"]}},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"TirUtilities.Vector3Extensions.IsZero(Vector3)","commentId":"M:TirUtilities.Vector3Extensions.IsZero(Vector3)","id":"IsZero(Vector3)","isEii":false,"isExtensionMethod":true,"parent":"TirUtilities.Vector3Extensions","langs":{"$type":"System.String[], mscorlib","$values":["csharp","vb"]},"name":"IsZero(Vector3)","nameWithType":"Vector3Extensions.IsZero(Vector3)","fullName":"TirUtilities.Vector3Extensions.IsZero(Vector3)","type":"Method","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"IsZero","path":"","startLine":5112,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["cs.temp.dll"]},"namespace":"TirUtilities","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public static bool IsZero(this Vector3 vector3)","parameters":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","id":"vector3","type":"Global.Vector3"}]},"return":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"System.Boolean"},"content.vb":"<ExtensionAttribute>\nPublic Shared Function IsZero(vector3 As Vector3) As Boolean"},"overload":"TirUtilities.Vector3Extensions.IsZero*","modifiers.csharp":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["public","static"]},"modifiers.vb":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["Public","Shared"]}},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"TirUtilities.Vector3Extensions.NotZero(Vector3)","commentId":"M:TirUtilities.Vector3Extensions.NotZero(Vector3)","id":"NotZero(Vector3)","isEii":false,"isExtensionMethod":true,"parent":"TirUtilities.Vector3Extensions","langs":{"$type":"System.String[], mscorlib","$values":["csharp","vb"]},"name":"NotZero(Vector3)","nameWithType":"Vector3Extensions.NotZero(Vector3)","fullName":"TirUtilities.Vector3Extensions.NotZero(Vector3)","type":"Method","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"NotZero","path":"","startLine":5113,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["cs.temp.dll"]},"namespace":"TirUtilities","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public static bool NotZero(this Vector3 vector3)","parameters":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","id":"vector3","type":"Global.Vector3"}]},"return":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"System.Boolean"},"content.vb":"<ExtensionAttribute>\nPublic Shared Function NotZero(vector3 As Vector3) As Boolean"},"overload":"TirUtilities.Vector3Extensions.NotZero*","modifiers.csharp":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["public","static"]},"modifiers.vb":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["Public","Shared"]}},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"TirUtilities.Vector3Extensions.Invariant(Vector3)","commentId":"M:TirUtilities.Vector3Extensions.Invariant(Vector3)","id":"Invariant(Vector3)","isEii":false,"isExtensionMethod":true,"parent":"TirUtilities.Vector3Extensions","langs":{"$type":"System.String[], mscorlib","$values":["csharp","vb"]},"name":"Invariant(Vector3)","nameWithType":"Vector3Extensions.Invariant(Vector3)","fullName":"TirUtilities.Vector3Extensions.Invariant(Vector3)","type":"Method","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"Invariant","path":"","startLine":5114,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["cs.temp.dll"]},"namespace":"TirUtilities","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public static bool Invariant(this Vector3 vector3)","parameters":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","id":"vector3","type":"Global.Vector3"}]},"return":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"System.Boolean"},"content.vb":"<ExtensionAttribute>\nPublic Shared Function Invariant(vector3 As Vector3) As Boolean"},"overload":"TirUtilities.Vector3Extensions.Invariant*","modifiers.csharp":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["public","static"]},"modifiers.vb":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["Public","Shared"]}},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"TirUtilities.Vector3Extensions.Abs(Vector3)","commentId":"M:TirUtilities.Vector3Extensions.Abs(Vector3)","id":"Abs(Vector3)","isEii":false,"isExtensionMethod":true,"parent":"TirUtilities.Vector3Extensions","langs":{"$type":"System.String[], mscorlib","$values":["csharp","vb"]},"name":"Abs(Vector3)","nameWithType":"Vector3Extensions.Abs(Vector3)","fullName":"TirUtilities.Vector3Extensions.Abs(Vector3)","type":"Method","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"Abs","path":"","startLine":5116,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["cs.temp.dll"]},"namespace":"TirUtilities","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public static Vector3 Abs(this Vector3 vec)","parameters":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","id":"vec","type":"Global.Vector3"}]},"return":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"Global.Vector3"},"content.vb":"<ExtensionAttribute>\nPublic Shared Function Abs(vec As Vector3) As Vector3"},"overload":"TirUtilities.Vector3Extensions.Abs*","modifiers.csharp":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["public","static"]},"modifiers.vb":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["Public","Shared"]}}]},"references":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"TirUtilities","commentId":"N:TirUtilities","name":"TirUtilities","nameWithType":"TirUtilities","fullName":"TirUtilities"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","commentId":"T:System.Object","parent":"System","isExternal":true,"name":"Object","nameWithType":"Object","fullName":"System.Object"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System","commentId":"N:System","isExternal":true,"name":"System","nameWithType":"System","fullName":"System"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"TirUtilities.Vector3Extensions.IsZero*","commentId":"Overload:TirUtilities.Vector3Extensions.IsZero","name":"IsZero","nameWithType":"Vector3Extensions.IsZero","fullName":"TirUtilities.Vector3Extensions.IsZero"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"Global.Vector3","isExternal":true,"name":"Vector3","nameWithType":"Vector3","fullName":"Vector3"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Boolean","commentId":"T:System.Boolean","parent":"System","isExternal":true,"name":"Boolean","nameWithType":"Boolean","fullName":"System.Boolean"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"TirUtilities.Vector3Extensions.NotZero*","commentId":"Overload:TirUtilities.Vector3Extensions.NotZero","name":"NotZero","nameWithType":"Vector3Extensions.NotZero","fullName":"TirUtilities.Vector3Extensions.NotZero"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"TirUtilities.Vector3Extensions.Invariant*","commentId":"Overload:TirUtilities.Vector3Extensions.Invariant","name":"Invariant","nameWithType":"Vector3Extensions.Invariant","fullName":"TirUtilities.Vector3Extensions.Invariant"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"TirUtilities.Vector3Extensions.Abs*","commentId":"Overload:TirUtilities.Vector3Extensions.Abs","name":"Abs","nameWithType":"Vector3Extensions.Abs","fullName":"TirUtilities.Vector3Extensions.Abs"}]},"shouldSkipMarkup":false,"_enableSearch":true,"_appFooter":"TirUtilities","_docfxVersion":"2.58.9.0","_appTitle":"TirUtilities","_systemKeys":{"$type":"System.String[], mscorlib","$values":["uid","isEii","isExtensionMethod","parent","children","href","langs","name","nameWithType","fullName","type","source","documentation","assemblies","namespace","summary","remarks","example","syntax","overridden","overload","exceptions","seealso","see","inheritance","derivedClasses","level","implements","inheritedMembers","extensionMethods","conceptual","platform","attributes","additionalNotes"]}}{   �?  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib"}	   �?   